module MEF_main(input clock,				// clock de 50 MHz nativo da placa
					 input new_data, 			// novo pacote de dados recebido
					 input [7:0] command,	// requisicao recebida
					 input [7:0] address,	// endereco do sensor
					 input [39:0] data_sensor, // informacoes do sensor
					 output [15:0] buffer_tx,	// novo pacote de envio
					 output reg send_data_tx,	// sinalizar que um novo pacote vai ser enviado para o tx
					 output reg inout_sensor);	// iniciar o sensor
		
	// Declaraçao dos estados 
	parameter IDLE = 3'b000, 
			  READ_DATA = 3'b001,
			  CONTROLLER_SENSOR = 3'b010,
			  PROCESS_DATA = 3'b011,	
			  SEND_DATA = 3'b100,
			  INCORRECT_DATA = 3'b101;
		
	reg [2:0] state = 0;
	reg [23:0] cont = 0;
	reg crt_decoder, // enable do decodificador para casos normais
		 loop = 0;	// avisar que esta em sensoriamento continuo
	reg [7:0] reg_command = 0;	// armazenamento do comando em execucao
	reg [7:0] reg_address = 0;	// armazenamento do endereco 
	reg command_invalid = 0;	// enable do decodificador para casos de erros
	reg [39:0] reg_data_sensor = 0;	// armazenamento dos dados do sensor (para nao perde-los ao reiniciar o sensor)

	// declaracao do modulo referente a tabela de comandos
	commands_table a(reg_command, crt_decoder, reg_data_sensor, command_invalid, buffer_tx);
	
	// verificacao do loop
	always @ (reg_command) begin
		if (reg_command == 3 || reg_command == 4) 
			loop <= 1;
		else 
			loop <= 0;
			
	end
	
	// armazenamento do comando atual
	always @(posedge clock) begin 
		if (loop) begin 
			if ((command == 5 || command == 6) && reg_address == address) begin
				reg_command <= command;
			end
				
		end
		
		else begin
			reg_command <= command;
			reg_address <= address;
		end
			
	end
		
	
	// maquina de estados
	always @( posedge clock) begin 
			
			case (state)
			
				IDLE: begin
				
					// Saida dos estados
					send_data_tx = 0; 	
					crt_decoder = 0;
					inout_sensor = 0;
					command_invalid = 0;

					// Transicao de estados
					if (new_data)
						state <= READ_DATA;	// caso um novo pacote chegue
					else 
						state <= IDLE;	
						
				end
				
				READ_DATA: begin
				
					// Saida dos estados
					send_data_tx = 0;
					crt_decoder = 0;
					inout_sensor = 0;
					command_invalid = 0;
				
					// Transicao de estados
					if (reg_command < 8'd7 && reg_address < 8'd32)
						state <= CONTROLLER_SENSOR;	// caso esteja com a info correta ou em loop
					
					else 
						state <= INCORRECT_DATA;
					
				end
		
				CONTROLLER_SENSOR: begin 
				
					// Saida dos estados
					send_data_tx = 0;
					crt_decoder = 0;
					inout_sensor = 1;
					
					// Transicao dos estados
					if (cont == 24'd12500000) begin	// temporizador referente ao recebimento dos dados do sensor				
						state <= PROCESS_DATA;
						cont <= 0;	// contadora zerada
						reg_data_sensor <= data_sensor;	// armazenamento dos dados do sensor
						
					end
					
					else begin	// persistencia no estado ate a contadora chegar ao final
						state <= CONTROLLER_SENSOR;
						cont = cont + 24'd1;		
					end
					
				end			
			
				PROCESS_DATA: begin
				
					// Saida dos estados
					send_data_tx = 0;
					crt_decoder = 1;
					inout_sensor = 0;
					command_invalid = 0;
					
					state <= SEND_DATA;
					
				end
					
				SEND_DATA: begin

					// Saida dos dados
					send_data_tx = 1;
					crt_decoder = 0;
					inout_sensor = 0;
					command_invalid = 0;
			
					if (loop)
						state <= READ_DATA;
						
					else 
						state <= IDLE;
		
				end
					
				INCORRECT_DATA: begin
				
					// Saida dos estados
					send_data_tx = 0;
					crt_decoder = 0;
					command_invalid = 1;
					inout_sensor = 0;
					
					state <= SEND_DATA;
				end
				
				default: state <= IDLE;
			
			endcase
			
		end
		
endmodule 


module commands_table(input [7:0] reg_command,
					input crt_decoder,
					input [39:0] data_sensor,
					input command_invalid,
					output reg [15:0] buffer_tx);
					
	// quando qualquer uma das tres entradas mudarem
	always @(reg_command, crt_decoder, data_sensor, command_invalid) begin
	
		if (crt_decoder) begin	
		
			case (reg_command)
			
				8'd0: begin 		
					// caso de erro
					if (data_sensor == 40'd1099511627775) begin 			
						buffer_tx[15:8] <= 8'h1F;
						buffer_tx[7:0] <= 8'hFF;							
					end
					// caso esteja correto
					else begin 							
						buffer_tx[15:8] <= 8'h07;
						buffer_tx[7:0] <= 8'hFF;							
					end	
					
				end
			
				8'd1: begin	
					if (data_sensor == 40'd1099511627775) begin 								
						buffer_tx[15:8] <= 8'h1F;						
						buffer_tx[7:0] <= 8'hFF;		
						
					end					
					
					else begin 								
						buffer_tx[15:8] <= 8'h09;
						buffer_tx[7:0] <= data_sensor[23:16];							
					end
					
				end
				
				8'd2: begin
					if (data_sensor == 40'd1099511627775) begin										
						buffer_tx[15:8] <= 8'h1F;
						buffer_tx[7:0] <= 8'hFF;										
					end
								
					else begin										
						buffer_tx[15:8] <= 8'h08;
						buffer_tx[7:0] <= data_sensor[39:32];										
					end
									
				end
				
				8'd3: begin
					 if (data_sensor == 40'd1099511627775) begin 		
						buffer_tx[15:8] <= 8'h1F;
						buffer_tx[7:0] <= 8'hFF;								
					end	
					
					else begin 
						buffer_tx[15:8] <= 8'h08;
						buffer_tx[7:0] <= data_sensor[23:16];
							
					end
								
				end
				
				8'd4: begin 
					if (data_sensor == 40'd1099511627775) begin 								
						buffer_tx[15:8] <= 8'h1F;
						buffer_tx[7:0] <= 8'hFF;								
					end
						
					else begin 								
						buffer_tx[15:8] <= 8'h09;
						buffer_tx[7:0] <= data_sensor[39:32];								
					end

				end
					
				8'd5: begin
					buffer_tx[15:8] <= 8'h0A;
					buffer_tx[7:0] <= 8'hFF;
					
				end
				
				8'd6: begin
					// forma inteligente (com uma linha so) -> buffer_tx = {8'h0B, 8'hFF};
					buffer_tx[15:8] <= 8'h0B;
					buffer_tx[7:0] <= 8'hFF;
					
				end
				
				default: buffer_tx[15:0] <= 8'd0;				
			
			endcase
		
		end	
		
		// Caso algum dado do novo pacote seja invalido
		else if (command_invalid) begin
		
			if (reg_command >= 8'd7)begin
				buffer_tx[15:8] <= 8'h0C;	// comando invalido
				buffer_tx[7:0] <= 8'hFF; 
			end
			
			// caso o endereco seja invalido
			else begin
				buffer_tx[15:8] <= 8'h0D;
				buffer_tx[7:0] <= 8'hFF;
			end
			
		end
		
		// caso nao seja nenhuma das duas opcoes
		else 
			buffer_tx[15:0] <= 8'd0;
							
	end		

endmodule